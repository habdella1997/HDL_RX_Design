`timescale 1ns / 1ps

module datagen #(
    parameter PHASES  = 16,
    parameter WIDTH   =  3 //QPSK -> 2 bits {-1,1} , 16-QAM 3 bits {-3,-1,1,3} , 64-QAM 4 bits {
)(
    input clk_i,
    input rst_i,
    input enable_i,
    input [1:0] modScheme_i, // {QPSK = 0, 16-QAM = 1 , 64-QAM 2}
    output [PHASES*WIDTH - 1 :0] data_o_i,
    output [PHASES*WIDTH - 1 :0] data_o_q
    );
    
    localparam integer PAYLOAD = $clog2(4096);
   
    
    
    reg [WIDTH-1:0] data_i_reg [0:PHASES-1];
    reg [WIDTH-1:0] data_q_reg [0:PHASES-1];
    reg [PAYLOAD-1:0] read_addr;
    
    integer i;
    always @(posedge clk_i)begin
        if(rst_i)begin
            read_addr <= {PAYLOAD{1'b0}};
        end else begin
            if(enable_i) begin
                read_addr <= (read_addr + PHASES >= 4096) ? {PAYLOAD{1'b0}}: read_addr + PHASES;
            end
            for(i=0; i<PHASES;i=i+1)begin
                data_i_reg[i] <= {data_ext_i_sym2[read_addr+i],data_ext_i_sym1[read_addr+i],i_data_sym1[read_addr+i]};
                data_q_reg[i] <= {data_ext_q_sym2[read_addr+i],data_ext_q_sym1[read_addr+i],q_data_sym1[read_addr+i]};
            end
        end
    end
    
    genvar j;
    generate
        for(j=0; j < PHASES; j=j+1)begin
            assign data_o_i[(j+1)*WIDTH -1 -: WIDTH] = (enable_i) ? data_i_reg[j]: {WIDTH{3'b000}};
            assign data_o_q[(j+1)*WIDTH -1 -: WIDTH] = (enable_i) ? data_q_reg[j]: {WIDTH{3'b000}};
        end
    endgenerate
    
    /*Scaling*/
    
     
    

    parameter i_data_sym1     = 4096'b1110011000100000011110000000001010000010001001110111000011110011010001111110110010101000011100101011110001111010101111100011110101010110100110111000000111010011011001111111000000010001010101011111010010001101000010111001110101100110100001100100001000010001111000111000111100110000010011011100011101010100011000101010111111110010111011001110110100100111111100000101011011110000100100111110010111110000100011011111010100111101111100100011101111101000111101000011010100001000011101011110011110100100001100110110011000111000110110110110011001110111100001111110010010100110101111100100001000101011010001110111000011011000110011011110011011010000110000100100101000101100101111010001000001010100001011110010000101010101101101100100110011010000100111111110011000110111110000110111111001111110000010111001100001101001000000101001011110110101111000110110001101100011011010110000111001010010011110011000111101001111001110101000110100100001000000010111010011010010011101010101000000000010001011110101101001000101000000110011001011011010100110111101100011010011100011001010000000000011000101111011000100101110001010100011101110100111001000000011101010110100101011101010100111101011110111001010110111001100101101101110100100110011001000010110101101001101110111111111100010100111101000110011001111001111101101001000011001100011000010001100100001001010010110001110010101010100101001100001110010111010101010000101001100011111111111001001010100001101001101100001100111110010010110100001110011101101110000111110011010011000100010001000100101011101101000001100010011011101001110101000011111000101111000011100010100100111011011111010011011010110001001101000001100100001010010001101000000111001001010001000101000000100010110010110110010010101101010111010101011000000001111110000100111111001111101010110010001110100011101011001000001011010011001001000100101001111100110111000001010110011111101001100000000011011010001110101001101111100001101100101110110001101011010011101100001001010001101010011110000010000001010010011101010100100001101100111011000011101010000110000111001100110011011100100000100010001111101010010100101000111100101110100011011010001100000101000111110011100000001111100001001111010101100011100001111101010111100010001010010001111100010101001111010000011100110110010100000001010010000110100001011110011001000011110100010011110101101110011101100100011011110100010101101010101110101010011000100001011011101111000000100011100000010010111010111001111110000011011011001011110000101000110111101101100100100100001001011100010010001000111010100010010100110001111011100111100000101111110011000011010011001100110010010110100111111010111000100101101010010110000101000101001011100100111010111111010010001110001111110110110010111000100011000000011110000000111101111011100000100101111101100001000001110011101100000001010000111010011011101001111001011010101001110111000111110101010001111101001101111110010110000110100001000001111000100000100011011111011000010101011011111110110011010101100011110001001011011111111101011000110011100101101001001110111101110001001111110000110000000000000011001110101100110101000101011000010000110100101100011111011101101001011100100110101000111010100010111110001001001101010011111110110011111000001101000101001011111100001111111001011011000111000001101010110111011000011001110011011000010010101010101010101011010001000000111010110101001100001011010000011110100000111110010000110001011001100110100101100111010000000110110011110011011011000100100111000011001000110010110101111010001111011011101000101101001010111011101001010001000100001011111111100110000100010011000011110001100100101010101010111011101001110010010000000111001111011100101000101100101100111100011000010001011111011001001000000111100011110001101001100000110110111111100101101010100100100100011000011001111010000111011100110110011100100011001000001101000011110111001000010000110110011001111100101111111000010100010000000111010000111111111100000011101001011101111100010110011010110010100010010011010110001111100000011000010011011011100000001101111000001010111000100110101100010000010001010011110000111101101100100000000010111;
    parameter q_data_sym1     = 4096'b0100000111010001111100011101011010101100101000001011010101001110010010111011011010011110001110010101100001011100010001000110100101101000011000011101101010011111011011101101000111111100001100000000111001011010010110111000011101110100011011000100101110110100001100001111110000011101001100011000100011100010000010111100111011110010111100011100101101001000101010101001011011111101010110011001001110001011111000110010101001010101001100100101010101110100011110011101000101100110010100000011000100001111100111000101100000100110000100010111001010101000010110011111010111110010011101110011010111010101011111111001110010111000100110011111100100010111110000000110000000101111000011100100011101100010101110101110101110000100010011100001011101011100110010111101110100101011010101110011001111000010101010101011011001001100011101011010110001111101010010010001011000000010110001001110110010101010100011100100101101000110001110111101101001001000110000111111000001100011000100010010111001011000001110001100100001111010110110010111100101001110101000001101011110110000110111011100010001100001101100100100000000010101010001111001001000011001101111101101101110101001001011010010100010001100101101000111101011111010011000100011110101000011001010011111101101010110101001100101011100000001100111111001000100111111101110100111111010101100001010010101111111101100111000101111100011010001100011010110000100001000110010001010111000101011110101001111110111000111001101010100010010011010101011111111001001110111001000000110000001000010001011110000000111100011111111001001010111100101100111110110100100001000000101001011001101000010001101110001000100010100011001111110100010011100000010100001011100101111000011011110010110101100100101110110101110111011000110000010001110001100000011001001010111110110010001100001111111010111000111011010110001011101110001101000001111010100110111011000011101011111111110100100110000001000101101011000010001010100111111101011100010010110000101010110100100011011101110010000010111110000110110011000000011100010001101010010110010000010100000110101111010011101001110101001111001010010010100111101100010101111100000000001010001100111100010101111010011000010011000101011111111000111000111000111001000101010010000000101100101110011011010101010100111000110100111111010101000100110100101101010001100110010011001011101010101101101111000010011010010101101110010011000000110110011100111010100101100111011010101010001100000011101111000110011111010000100101011011010011011000010100100100000010100110111001111000110010001011100011111110010110111001111011010110001110000000001010001010111110111101000111000001011000011000110100111000100010101011110101011000000110001010111010010100010010011000110101111000011000100100001101101010010001001110100110110011010110110111111110101000000011011101110000001100110110100000001100000011010011111000100110010101110100100110000011001111000001100100000110100100101101000001101111000001111010000000000111001111000010011111101000111011000111111010111100011001111100101011011000001001000011011011111010010111111111111110001101001110010110000100100010101111101110010000101111000111011110110101101000100110001111011100000110101111100010011101001100001101000011011010000100001111100011111001100100011011101011111011101100101000011100111111111000110011011101011111100000111001100101001110000101100000010101101101110010111011001110011110101011101011001000111110010010110011101011001011011101011111011111101100101001001110101100100000011110110100001111000001110010001001001011010011110111011000101000011001010110100101001001010010001001010101111111010110100011100111000100110010101111111010010111010100001111011010010010000010111101011010110111101011000010100010010000111001100010101011100010011000101011111000011001100111101101100011001101100010111011000011110011000100011001000101000100110111001011010011011111000101010100100110011101111111110011000001011100100011001010011110011010110010110001110000010101100100010100010010010100110001011111111001001110100100111100011010111110100011110100000001100110101111100010010011011101010000001110111101010100100001111101010110001101111010101;   
    parameter data_ext_i_sym1 = 4096'b1001010101010000000111110010010010111010101001001101111001011111000001110011111110000000001000000010100110111000101100111000000110101101111000111100100111000001010001100101100010101001011100010010100110010001011010001110000011000001011010100011011000010101000001111000000110010100001100000101110110110011000100111100010010011101101000010101100001101001000010110010110101110100101100011101100100101110111100001101000100000011001000111110011101111001100001010111000100101100111011001001000000100111010011100100101100011001000101110101100111011101100010111111001001101010101010010000011001000111001000010001001011010001000000001111000000100100000111001110101101101001000101011100101101110111011000000101010100111011010011001111010111001100100110001010001110111011001110110000110011101110011010001001101100010110111110110011010101111000110010000000000000110110010010010110011010110101010010111111011000011111001011011010001100110110110111101111100000100001010011100100001110110000111111101100010100011111111010110101010101110000111000011010111110010011010111010100001110110100010101001011011011010110010101001010110110101010011110010001011001110100111010000110010011000011010101101110100001101110101101001110110111110100001000110100011110011011100110000001001011011110000100011011010001000111010110110010111010111111101000100101111010111001111101010111011100111100100101000010101110100100110010100000001011001110110010010001100110010001011111100100000010110011110000101100101100101011011000101001011111111110111111111110010100100001001011110000100011001100001100010110000000111011111001001000110100001000110010101110111110111011010100001001100001111110000101000000100001011000001011011110001100101111101101000011111011110001110010100000000000100001010111010100101001011101100010110011010111100011111010010000101000000110011110010000000001010110000010010100101011011101110110011101101110100000101110001001100110101110000110101101001111100110101011101100010010100101001100100111010101000010011110100001010111110100101000101110010010001101001110110110101111100011100001010101100100010011010010100101101111001101000010110001110000110010010100100111110100110110001011010001001000101100000001110011001100011111110001011000111000101111101100010011100110011001100100000111011111110110110110000011011110010110100100110000001011111110111010101110000000101100100100010111010000110100100100000001000111000011011101010000000000101001001011011100111001100111101001101001000010101100010111011111110000111110000110001011111100011000001001011011010001100110111001010110101111110111011110110110101000010011101010110101110000110010110011011001101110001101111001111010001110000101110110110001000100001000010110100110100110101010010100000001000110010110011011011110010011000110010110000100000111001000010011010111110011101110010001101011101000010100001011101111110011110000101011111011001001011111011000001000001110101000010011110001010101101000110011010110001100000011001010111100010010111100011011011010000101101100100011001101000101000100010010101001111001101110100011101111111011111100100001010000000100000010001101100111010011010011110110001001000010000001111111011010100111101111001000100000001100010101011111100110000101101100001110000001110000011111001101111011011000110101000000111100111101010101100101100001000110001110000011000001110100000100100101010111100111111101111000011111101110110100010011110101101000000011101100100111011010110110000011001000000100010100111001101101011011111000011111001011000110101100111110100111100001011011011011101110101111010000100010111010010011001101101100111110000100101100011111100110111001110000100101010110000100011010111100101010010011010100111110100011101111101110000111101111101001011101101011100101011111110100110000110100100100100100111101001001101001010000110000110000100111011011001001111000110100011011100011000111010001001010001001101010101001111100100101010111010000010011010110101000000010110100010001001110100000001011100111101110000001010101111101100110000000111000001110001100111011000110110111011100101101000010010000100111110000011101001000010010101101010111;           
    parameter data_ext_q_sym1 = 4096'b1110001100001101000000110110010000110001011110011011001001001010110101001011000000100110111100000100011110001101101111000010000000011011000010100001111100111101111001110101001101110100101000000101000001111000110111011011001001001110110100001010100000011010000110111010101001110011100101100010101111011001010000001111101110011011101111001111111010001101001001100000101001010011011000011011100000110110110001111011100000000110011000101110001101011100010100010111111001000100101101111111110000011010010001001000101000100100111100001111011101001000111010111000001100111001110100010101100100100111100000011000001010111100110000010110001101100100001111001110000001011001010101010111010001110001101101111001110000110011110001000001101000010010011110111000010000110100110100100111011000000000001111110010001110011011010010101001001001011111100100110100011100100000010010001011100110101111111100101011111011011011110010111110111101101101001110011010001011101010001011111001001111110110100011011101011110110010001000111110111111001111110100110110111110100000111101100010101001011111001000110100111010011110001101000101111111111010011111101100110100111100011111010011011011000101010110101011101010110010010111110001100110101001011100111100000100000101010010011010000110110100010100101100100111111101111100011010000000101100111111100101100110100000000000010110011011110101001110010100011001001111110100110001100101110101101110000010110010110010101000000110000111010111011001010110011111110101110100111010110101001101000101000001010101100011001100110000000001000100011001011111111000010010111110000111100001000011010010100101111011101011001001011100011100011100100011101100110100000001110010001111101011010000011010000010101100000001111110000100011100101111111011111010010001111101011101000011101000001100001010101100100001010011011010111100101000111100000010010111100100000110011110101110010011100000000110000100100101100101100111001111100101001001010101010101010001001111010000110111011111011001111010111100011100101110100000111011101110111010110110101000100010100000010110100001000101101011001000010000100001010111101111000000010101000100001110101010101110100010011111100010010100010000011011000000011011001011011011010000000001001100100100001000101001100001001111010000111000101000100111111100111001010001010111110100011011100001100010000011111000100111110000001000111111011100000100010101101110110001100101110011111101100001110111011001000010111011111101100110010000110101111011001001101100010111000101001011000001101010010000000110100101111010010000000011001100010110101000110110011011011111100001110111111100001110001010010001000001000000011000011001101011001000000001101111111000010010101001100110011100011110010001110110011101101001111000110000101110001110001101001111100101011100011010000111110001111000000110000111110101000110100111011111010011111100011100111110011000001001100011011111001011111100100000010010001111111100001001000101010100110000111010111101011111110100010101110111101011110100101011010000100001100101100000001100010010001101010101101010001001101111001110110101101011001001110110001001001111111000101111001101111001100010110011010000011000111100001001010110010101010000100000001101100011011010000000111110000101011110110001000100001110110011110101100110001110101110010000101010011100110111010110001000111001011100001101010011101101000111000001001111111000010100000000111000111111000111011101100101000111000111110100111111101101010100010100001000000000110010001110111101001010100011101011011110011100111100111101010101110110001100110110010100011101110100001111100011010001000100001101001011010101010001011100011000011101001010100110101011000101000000001000010101001010010100001101101011010000011010001010100000110010001000001010111011101100010111011111100000100111101111101000111100010100100001110001111101011000001010110001000001011001110010001111101001100101011000010101011011011010000010001011100000100001011001010000010110110010110011011001101000011101000101011111000001001011011010010110100001011101101001010101011011110010101001001101101001111001001110100000001100101100111100;     
    parameter data_ext_i_sym2 = 4096'b0111000111011000010010000101101001110010000101011011111100000010010101100111100011000011100111101000010110010000111110111100001101000010110110000011001000101101011101000110101010100011011110011100111110011001001110100111110000101111100100101110010111001001111011011111001111111111100010010100100110100111111010000111000011101111000100001100000001100111100101110101101100000100101001111100111001011011011101001001111000111100010100011001011001001111001101000000011110010101011101111101110011010000101111011011111011000110101110000111111110001101100111111110001110000100101101110100010010000001001010000000000011011011001100001001001111001000000001111001110000110110000000010101001110011110100010010100100001010111000111011001110100011101010000110101110110011111000101110101001001111100011001011101111110110111001101111000100011001000000010110101000111010100001010100100110010001100010010100011101001000001011000101010011010110001100111000101011100011111010010010100001010111000100101001010011101001010011111110001101101101011101101010001010011011100101111101001111001000000001001011001101010111100001001111001101001110100111111000010001010011011011111111111011010010111001110111011101101100101010111101000011001000110011010010100101000101010111111001110001000010100000010111000010011100100000011100011010111110101110111000010100110110111010000111000101101011001101110110010100101010010101010000101001100011011110000110001010011011101010001011010101111011101110101011010111110011110101000010000001110011000001111111000110101000000110110000101101010110111110010110010101010101100011100101010011100110001000001010111100111110011010100101110001111110101110000011000111011010101111000010111011011010000001110010010110010010110000010111101100100001110000010100011100101000010000111101001010111110101110010001100011000110001011000111101101111110010000110001101111010111101110001101111110111110000110010111001101010100001100111001010101010111111010000111100000011111011001011000001010100110100001001101011100000100101000010100101111000110101011000001110110110000111001101100100001101110011000110011011010111101101101101000110010111101110100011110101111001000100110000011101011010100101011100001111110111000110100011010111011010101100000100101111100010111101100111111000111011110100011111100000001000100100000011101001001101100000111011101000110000001000111010111110101000001001011110100101111001011100001000110000110010100011000000100101011110100010111100000001101001001111100001011111010101100101100010101110111100101101011100111000100101110011101111110000000011011001110000001101000111010110110101111101000010100100101001000010110101010011001111110011001100000010110101011001101010100001010000000011001110111100110000110000111011100000001001111110000011101101001001100010011011001010000001111010111110010110111111100101101100001010011000010001101001111010101001010000101101110011101000100100011011011101100001001010000011011100011001111011011011100101101101111011110100011111100011001011001111011101100100011101111010100010100100100011110010000101010011000000001110010011100101110011100111011100100101011000011000101110100110000000111011111101111001110011101010011010000100101010000011110000110011011001110011011111010101000011100001000011000001110011101011101000100101001001110011111001001100011001011010010110000000111001001110111111011100111111111001000000110010111010110001010111100100000101010110111101001011110000001101001110111111111010011101011111100110101111001101011001111111000101110000011110110101101110100011110000000000111001000000100100100001101101000001000111110111100010010100010010110101010100001011100100111010010001111000001000010010001110100001111100101000001010001010101110001110001110110111100101111000000110010001010100111111100010011101000001011000100011011111110001101001001101100101110100001001010110001000001001100010111000011110001110010111000001100001000110111011111011101101110010101010000110101110101011101010010000110000110001100110001001010010110101010011001100010010000010111000001000101011000011110010100101111110010001101111101011001010011101111100101011000110100100;
    parameter data_ext_q_sym2 = 4096'b0000101001101111001010010111111100001110101100011100110010001111101010000001011111000110010111110110000110010011000110110010011111010011010001101010010011000101100001001010111100110000010011110110110000010111100111010110100111101101010001001100001110111111011101100111010000000010010100111110000110110000010011100100110000000111000001110100011011000101010111101001011010001111001000110011010011011111000011000010110001101100111110111000001101000100010111100101111110100100011101100011101111001110100110000110111010000000110111011101110011010111101011101001010011011101110111011001011100101000110001011101001100101100011011010000001110001100100110010000010011110101011011101000010100000010001100010000010100101101010101111110000010100111101000001100001010101010011111000100110000011101001001010100100000010000101011111001001011110000110010001111001011111100010101011001001110011100000010111011111101010011001010110001110000111011110010011100111111011101010100010010111010001011001110000010011010001000100001100000111111010010010011100111001010111011011110001110010010000100010100011011010111101001110110000111101010100101010000000011011010101100101111110001101001010110110010000100001010010110010000100100101101001101111001010001010001000011011011001100011101100110101111101000010110100100110111011110000101100110011010000000001001101110101101010001000110000010001110000111101001000110100111011101100011111000001000011101110111101010001011000110011110000000111101010100101111101110111000110000110101000111000101110001100110100111010010110000110011001001111100001111001111110110101010100010011101001110001000101010110101100000001001000110111110001111011111010110100011101100011101001010101001011001111101100001000110011000011010110010011010111011000010010101110100010100101011001100110001010011101100001011110001010001101011010101011111000101100000011000110011010011010101101110110100111010001111010001110010110110101111010110011000101010101011011000110111111010001100010100001000000110010000101001010101010101000001101101110100011110000110000111000110101111000011010000000100010111100010010110001111100100101101000000001100001100010110111001111110111101100000011110010111100101011100101111011010001011001010010000110110011110111000100001110100000111000111010111101100000100111011001111110001110100111000011101010011001000011110000011011111111001001011100111001010000110101011111111101010100010011000100001000001111101111011100010010101111000110101100011000110110011000100110010010110011110100001000110001111011001101100010011000110111100111011001101001111010000000010011101000100011011101010001010111110101100011111001110000010101000110010011001001101101001000011100000111010011000101000101111111000001001000001100010010001110111010010101110010110001000100111001011011010001110101000101000110001011001100000010001100100000110100110011100001001001110110010100010111110110010100100101110011110000010001111010011001000010011000111111001001011010011101010100011100010111111010000001010111101001011000110011001001100001011001110111011000001001001111010101110011011011001101110100001010011010011011011101011011100101000010001011111100011101000010011101101001101110101001000101000000110010011100101101110000100010001011010110001010101010001010111000011101010001100010111011011000101110100101000111001001011000110011000110100010100010100000011000001000010010110101001111000001000111010110010100000010111000110010111001100111100110010011101111000011110000011001011101010011111011110100101001111100011011001110100101011010100001000011011011110110101100100000001100100011111010111001110111111110011100110010101110100111000111100000101011101100011100101101010100101010100010110100111000111000001110010100101100110100000100011000000010111000101101000010011011000111000011000000000010100001011111010001101000001100110011001010100101000100011001011101110001100011000111010101111001000100001110110111100100110111000000010110110101010101101010110001011010010010110010010100011100001101010000100111011000000111101101111000111001100110011001001010100011011101001100110100100110110100110000001001100100100000100011010;

endmodule
